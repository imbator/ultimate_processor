module mux(
);
endmodule